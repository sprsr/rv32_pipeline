module rv32(

)
