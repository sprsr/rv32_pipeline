module debug_port(
    input [31:0] registers [31:0],
    output [31:0] reg0,
    output [31:0] reg1,
    output [31:0] reg2,
    output [31:0] reg3,
    output [31:0] reg4,
    output [31:0] reg5,
    output [31:0] reg6,
    output [31:0] reg7,
    output [31:0] reg8,
    output [31:0] reg9,
    output [31:0] reg10,
    output [31:0] reg11,
    output [31:0] reg22,
    output [31:0] reg23,
    output [31:0] reg24,
    output [31:0] reg25,
    output [31:0] reg26,
    output [31:0] reg27,
    output [31:0] reg28,
    output [31:0] reg29,
    output [31:0] reg30,
    output [31:0] reg31
);

assign reg_1 = registers[1];
assign reg_2 = registers[2];
assign reg_3 = registers[3];
assign reg_4 = registers[4];
assign reg_5 = registers[5];
assign reg_6 = registers[6];
assign reg_7 = registers[7];
assign reg_8 = registers[8];
assign reg_9 = registers[9];
assign reg_10 = registers[10];
assign reg_11 = registers[11];
assign reg_12 = registers[12];
assign reg_13 = registers[13];
assign reg_14 = registers[14];
assign reg_15 = registers[15];
assign reg_16 = registers[16];
assign reg_17 = registers[17];
assign reg_18 = registers[18];
assign reg_19 = registers[19];
assign reg_20 = registers[20];
assign reg_21 = registers[21];
assign reg_22 = registers[22];
assign reg_23 = registers[23];
assign reg_24 = registers[24];
assign reg_25 = registers[25];
assign reg_26 = registers[26];
assign reg_27 = registers[27];
assign reg_28 = registers[28];
assign reg_29 = registers[29];
assign reg_30 = registers[30];
assign reg_31 = registers[31];
endmodule
