module wb_ctl(
    input
)
