module branch_comp(
    input [31:0] i_dataA;
    input [31:0] i_dataB;

)
