module instr_mgr(
    input        clk,
    input        rst,
    input [31:0] instr_de,
    input [31:0] instr_exe,
    input [31:0] instr_acc,
    output       stall,
    output       hazard,
    output[31:0] data_a_mgr,
    output[31:0] data_b_mgr
);

reg [3:0] r_conflict_map;
reg [2:0] r_wb_acc;
reg [2:0] r_wb_exe;
reg [31:0] r_data_mgr;
reg [31:0] r_data_a_mgr;
reg [31:0] r_data_a_mgr;

//Function checking if the instruction is a write back instruction
function [2:0] write_back_check;
    input [31:0] instruction;
    case (instruction[6:0])
        // LUI Instruction: 
        7'b0110111: begin
            write_back_check  <= 2'b01;
        end
        // AUIPC Instruction: 
        7'b0010111: begin
            write_back_check  <= 2'b01;
        end
        // JALR Instruction:
        7'b1100111: begin
            write_back_check  <= 2'b10;
        end
        7'b1100011: begin
            write_back_check  <= 2'bx;
        end
        7'b0000011: begin
            write_back_check  <= 2'b0;
        end
        7'b0100011: begin
            write_back_check  <= 2'b0;
        end
        7'b0010011: begin
            write_back_check  <= 2'b1;
        end
        7'b0110011: begin
            write_back_check  <= 2'b1;
        end
        default: begin
            write_back_check  <= 2'b11;
        end
    endcase
endfunction

always @(posedge clk or posedge rst) begin
    if (rst) begin
        r_conflict_map = 4'b0;
        r_stall = 1'b0;
    end else begin
        if (instr_acc[11:7] == instr_de[19:15]) begin
            r_conflict_map[3] = 1'b1;
        end else if (instr_acc[11:7] == instr_de[24:20]) begin
            r_conflict_map[2] = 1'b1;
        end else if (instr_exe[11:7] == instr_de[19:15]) begin
            r_conflict_map[1] = 1'b1;
        end else if(instr_exe[11:7] == instr_de[24:20]) begin
            r_conflict_map[0] = 1'b1;
        end
        if (r_conflict_map[1] || r_conflict_map[0]) begin
            r_wb_exe = write_back_check(instr_exe);
            case (r_wb_exe)
                3'b00: begin
                    r_stall = 1'b1;
                    r_data_mgr = 32'hx;
                end
                3'b01: begin
                    r_data_mgr = alu_out_exe;
                end
                3'b10: begin
                    r_data_mgr = pc_4_exe;
                end
                default: begin
                    r_data_mgr = 32'hx;
                end
            endcase
            if (r_conflict_map[1]) begin
                r_data_a_mgr = r_data_mgr;
            end else if (r_conflict_map[0]) begin
                r_data_b_mgr = r_data_mgr;
            end
        end 
        if (r_conflict_map[3] || r_conflict_map[2]) begin
            r_wb_acc = write_back_check(instr_acc);
            case (r_wb_acc)
                3'b00: begin
                    r_data_mgr = dmem_out_acc;
                end
                3'b01: begin
                    r_data_mgr = alu_out_acc;
                end
                3'b10: begin
                    r_data_mgr = pc_4_acc;
                end
                default: begin
                    r_data_mgr = 32'hx;
                end
            endcase
            if (r_conflict_map[3] && !r_conflict_map[1]) begin
                r_data_a_mgr = r_data_mgr;
            end else if (r_conflict_map[2] && !r_conflict_map[0]) begin
                r_data_b_mgr = r_data_mgr;
            end
        end
    end
end

endmodule
