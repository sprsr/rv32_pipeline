module execute_ctl(
    input clk,
    input rst,
    input [31:0] instruction,
    output [31:0] instr_acc
);
